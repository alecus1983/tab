BZh91AY&SYD��U  �߀Ryc����߰����`>-�^��n �a����(m�����Ayڍ+�)�u� yǻT� $�FB����)�C�42�چ� 4Hʒ��4��    4�#��i�`��244@�I��=ML�4���A���ML��2e6�b)�����z�����2�M4��(���F�  4�⨤�Q!�� �E�UK	��� �� ��|�~���?����r��/��RPS���ànƄ�Lc�T��i�T�bI&��4�QD���D�`��N����io��1�i�/#��^\P������5@6@��>���|Zx��/��ssO�w��Ͱ��l�Z�� p�TY�f2�3��:x�(e#I'�-��Դ��o�X��|���1�84�����S�P��/������5\:c$��fӶܐsC�zm�Փf��)��+�0������"Sى��Ed�ו��}��i�;x<S�'	���4�p5�[�X��Ŗ]��L�fta/�L��X��7(�2�8�:�h=�ԏ��t�>�0�JP�l���*�����V�1����i�*K)�ܡ��1sFI9�z5'*N���ُ�8^�V�ub,��M
J[/P�%^�?o6�g���=t������Xȴ(fZ��pw,������ew�K	���jl��&�8�)�ʇuD��f4U��B,ZLda��H���b�8�cYH2Ca�K��8ދUk̄en�:�"l�cWpvXR*���[�l�8��!d)���6��V�:MkZ��J��!A�=�b���D�T���j�⡘�jT��u�L�p�Q�^0�)r
a�^��j�r����ʯ����o7/��kvv}|��L�^:4Zb����"�PL��N��h�"�3�
@�5�N�.�P?+�����xM��ُ���8�l_S���$D��x$!�*0*��A�$C���	�z�C6��4���i�87~Ǜ�z3\�'�Mk�E�`@!7�#�SU2���h8�/jX@���[`��O���{ �5Xu�ڶ�;�X�>8�8����MjWTãc6�cSe��5�c�er2R��� �3� D㓗�I��6Ӭ��#�`�����hps�/���c�S�s��� U��=i��m�n<[�0���чvQ�C�sƬ&:롪NɢFh��yIU�q�$^ք�q
��>O~���{q�A��~,�;Z�X�MC�H�ħ�Gr\fN9�6b�e3���6OR��}l��E�[4D�E�2c��>�+!¯�Y��ѤN��G��2��Q��F������t��d����n2�����L��c��a�*&�\��2������&fd�KA,L�`��1�+�$u�fR�NE��1F�Y� �;��0�T�g��<�<4Dd��L��ƭ�u5KJki@��A�li�G���j�7�V̚�y������>A�Z���UQ�oK��1A����O�$��i�����k��Fy��Zֽx�s8o
����r�'<u��n9�%��44��%�$���Y�U��l��-��.�$�8bs��-9��g���3Ժu�ɦ8�TV���b}�BGg��qǲSF;�x��6��H���,�㖮�M�9�:v��d=x9�R8�9:��Y�%�R��K�]��+)a�O��xOQ�fQD�n2�'n�|TX�y���{|��6�#�1G2�k��Jpi�z��%K�:���զL�Z�a���0�,ru\�9�����tm�hǔ�<p��mr��ă�R����9��=J��f���o�A?H��!����G:)�b�d��e�1U�&�ۤ��Q��4�S+��UC1���vT�i�KcS(���g��1�+}��0�5�sp�O2ǆ2a���b��/hp��
�l�۵S��,���6�#��Ԟ�o-���1�)uPF�NAI�Z�ptg_R���hF���Y]~L6B�4���`�G�*@�����hs�����,{P�#iz:�d~zA�:!!)�5d��q{��ꝲq�6߭u�h>��q㛮M*"����YlҸo�	�=����Qc"��J�S�a���+���ƭ�'�yQ=�4y�®�c�C��9�5YqƜ�O���/o)DVaj���kMۼ4m�����W�%���(=��S���c���C�F�U��R���5Uf�Y:��&c)HG)��Y��]2oILmx^>E�s'�-���,z�1I&Ni1�W�c+������D0������d:��������xRź���ǻ�*ԧ:�iA<s9>�i��2�SZBaԢ��GZ�:��T��YR��K^=@�w��f����o��|i�	�հ���H��;�KbhM���āP�ۉ��B��4�A��U�HL��Ļ��3�.����K��/�8���!@r��"+e�ޅ�B��w��C��V'P�f� $��:�Ne-��F�4_y2���HU:̋!y�k$|�+-�r�ͯ>��݁�P9j+N���1�K�S͍�$��5Pr�4m*%�h�\9�IE5�9�)*V�+�Leə�����>��Fv<��8i��d�'��6�A���#��V�+�*t��d��<�?��NQ�8�f-�HìI����'C�鬸VF�>ը��o��(ŉ�(��z���g�!���mQ�H���TKL��	�D3¶`�o�g��j�Ri�p�xr��1gr��/���mT�\�?�����EǓ�H��A��mB�8��.&�VUnj*mQtV��;�*��rNQ����N(r]B��W���=4���=��R�MèHiv%J��sT�_Ma���l��u���Q�&^�T�boL-5:�Cj�����z��l5ݙ��1�7�?�_��*o�.���Ar:�Ie*�PW�TQFth�ع�`ś��w������{# C�TA���HHH�"X�������@0�,��H�p�^��D����\U���C,J5�IF�h�M@j �
"�`���7B��@U��(�Ē�V@P��P�+e(��*!iDSf(���66�lϕ��lqK����07�Smܞ<-���b����ꦺ��W�Fo���~� �	X��Q��A�(�)~�M�X)����	!#�C�h��
�H�a �ax �E��#�������Ҿ�4��Z���
B��D���)�mWB�1�K4�o���V
�P�Ңq�z�ֻ�J4'L'Fh
7BH��[R,�5��B���О�}� �'GlBE�[�MAݓ�o7P�����P|Zx������������!בd�u�%��w�❣����!��$�u����}���8
�ep���F|�
�`���'�E����̡EB5*B�����)�>����u4��w�:|C��#����P��<�=��1_�q���6s���4ӽ�k\"�۴��oy���kC;�s��Cѵ^�z��L]��=��9>.w�����g[O�eϳ)��Ɋxp�2���>�l,������%"�) ���Tò�@[`���@�"ju�:�J�G� ���T��;Mw��PI]S#�{ԛH�ņ��3�D�}��ً3�qؘ�J�z��u�LV �	TGg>e�va���" "`�`1���88��m����ǁs�l8X(q/H{7���BCu�=����˭�!���l1��qlD7=�-��)t>�:�:F<��N}K�1v��4�(i]�֊�j�Q� �/�nCK^m�.Wg������p@���l��p�
%��3$EA<������b�����z�}�Аa|��:�����#G!̯pz�09�s���5?;(����Ǡ�Y_Ǌ�x��1W��u���{�ce��,��FR2є�Z�Nޫ4e������1tSJj����4`�[#�����6�lt0�=�t4�h��x���Q&�AEQ��Q��M,��
��p:��3�pp3��H'���
�X��3��v�0�C���x$�ht�3���� [ihP��牯%C$ԙ7XeGbEm���hp�;���D�ehr�"xa���#Ї~�Sa��Qz>��zPH?I��#��:�N�jݬ��3!<����,Bw��° �.-�W���dv:l;tކqjM�z��O:'051�G��hi�^-�?kH�&����؆��N�E���tH<�JE��C3����z~g��u=�d���	];���<�И��!�Il��l1��t��g^�8���Nt�ry1й����<���2E�!����᥁��φa���Ɵ�Ö��Ǔ��[�Pt���vn�6"nCpꥲ�4)���C�F�7�����#w: ru1�����o{�N�A` �ӭ�\���?� �=Z���V��1~;���h{�'V�L��pH��:hxp�4�g8f�6΅�}-{�h��`�}_�w�]��BA�IT